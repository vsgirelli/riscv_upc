package config_pkg;

  parameter integer ARCH_LEN = 32;
  parameter integer INST_LEN = 32;
  parameter integer REG_FILE_LEN = 32;

endpackage
